`ifdef 
`else
`define 
`include define.v

module (
	input wire;
	input wire ;
	output reg ;
	)

	always @(*) begin
	end

endmodule
`endif