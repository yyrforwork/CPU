`timescale 1ns / 1ps

`ifdef _REG_FILE_
`else
`define _REG_FILE_
`include "define.v"

module REG_File(
        
    );

endmodule

`endif